`ifndef MY_ENV__SV
`define MY_ENV__SV

`include "my_monitor.sv"
`include "my_agent.sv"
`include "my_model.sv"
`include "my_scoreboard.sv"

class my_env extends uvm_env;

	my_agent  i_agt;
   	my_agent  o_agt;
	my_model  mdl;
	my_scoreboard scb;

   	uvm_tlm_analysis_fifo #(my_transaction) o_agt_scb_fifo;
   	uvm_tlm_analysis_fifo #(my_transaction) i_agt_mdl_fifo;
   	uvm_tlm_analysis_fifo #(my_transaction) mdl_scb_fifo;

	function new(string name = "my_env", uvm_component parent);
      	super.new(name, parent);
   	endfunction

   	virtual function void build_phase(uvm_phase phase);
		`uvm_info("my_env", "build_phase is called", UVM_LOW);
      	super.build_phase(phase);
      	i_agt = my_agent::type_id::create("i_agt", this);
      	o_agt = my_agent::type_id::create("o_agt", this);
      	i_agt.is_active = UVM_ACTIVE;
      	o_agt.is_active = UVM_PASSIVE; 
		mdl = my_model::type_id::create("mdl", this);
		scb = my_scoreboard::type_id::create("scb", this);
      	o_agt_scb_fifo = new("o_agt_scb_fifo", this);
      	i_agt_mdl_fifo = new("i_agt_mdl_fifo", this);
      	mdl_scb_fifo   = new("mdl_scb_fifo", this);
	endfunction

	extern virtual function void connect_phase(uvm_phase phase);
   	`uvm_component_utils(my_env)
endclass

	function void my_env::connect_phase(uvm_phase phase);
   		super.connect_phase(phase);
   		i_agt.ap.connect(i_agt_mdl_fifo.analysis_export);
   		mdl.port.connect(i_agt_mdl_fifo.blocking_get_export);
   		mdl.ap.connect(mdl_scb_fifo.analysis_export);
   		scb.exp_port.connect(mdl_scb_fifo.blocking_get_export);
   		o_agt.ap.connect(o_agt_scb_fifo.analysis_export);
   		scb.act_port.connect(o_agt_scb_fifo.blocking_get_export);	
	endfunction


`endif
