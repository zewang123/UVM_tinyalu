`ifndef ALU_OR__SV
`define ALU_OR__SV
class or_sequence extends uvm_sequence #(my_transaction);
   my_transaction m_trans;

   function  new(string name= "or_sequence");
      super.new(name);
   endfunction 
   
   virtual task body();
      if(starting_phase != null) 
         starting_phase.raise_objection(this);
      repeat (10) begin
         `uvm_do_with(m_trans, {m_trans.op == 3'b011;})
		 `uvm_info("alu_or_rand_test", "op = 3'b011 , or_rand:", UVM_LOW);
      end
      #100;
      if(starting_phase != null) 
         starting_phase.drop_objection(this);
   endtask

   `uvm_object_utils(or_sequence)
endclass


class alu_or_rand_test extends base_test;

   function new(string name = "alu_or_rand_test", uvm_component parent = null);
      super.new(name,parent);
   endfunction 
   extern virtual function void build_phase(uvm_phase phase); 
   `uvm_component_utils(alu_or_rand_test)
endclass


function void alu_or_rand_test::build_phase(uvm_phase phase);
   super.build_phase(phase);

   uvm_config_db#(uvm_object_wrapper)::set(this, 
                                           "env.i_agt.sqr.main_phase", 
                                           "default_sequence", 
                                           or_sequence::type_id::get());
endfunction

`endif
