`include "my_driver.sv"
`include "my_if.sv"
`include "my_transaction.sv"
`include "my_env.sv"
`include "my_monitor.sv"
`include "my_agent.sv"
`include "my_model.sv"
`include "my_scoreboard.sv"
`include "my_sequencer.sv"
`include "my_sequence.sv"
`include "base_test.sv"
`include "my_case0.sv"	
`include "my_case1.sv"

